`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
//Ben Alexander
//Ryan Holland
//Ryan Zagala
////////////////////////////////////////////////////////////////////////////////
module mux(a, b, sel, y);
    input [31:0] a, b;
    input sel;
    output [31:0] y;
	assign y = sel ? a : b;
endmodule